
// SPDX-License-Identifier: MPL-2.0

`ifndef __OCLIB_LIBRARIES_VH
  `define __OCLIB_LIBRARIES_VH

  `ifdef OC_LIBRARY_ULTRASCALE_PLUS
    `define OC_LIBRARY_XILINX
  `endif

`endif //  `ifndef __OCLIB_LIBRARIES_VH
