
// SPDX-License-Identifier: MPL-2.0

`ifndef __OCSIM_PKG
`define __OCSIM_PKG

package ocsim_pkg;

  localparam DataTypeZero = 0;
  localparam DataTypeOne = 1;
  localparam DataTypeRandom = 2;

endpackage // ocsim_pkg


`endif // __OCSIM_PKG
